`define ADDR_WIDTH 9
`define DATA_WIDTH 32
`define STRB_WIDTH `DATA_WIDTH/8
`define DEPTH 256
